module sub_3();
	    implement code
endmodule
