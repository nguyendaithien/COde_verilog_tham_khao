module sub_2();
	    implement code
endmodule
