module sub_8();
	    implement code
endmodule
