module sub_1();
	    implement code
endmodule
