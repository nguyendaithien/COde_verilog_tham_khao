module sub_4();
	    implement code
endmodule
