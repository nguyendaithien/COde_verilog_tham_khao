module count_down( clk, max_sec_i, sec_count_o, min_count_o);
input 
