module sub_6();
	    implement code
endmodule
