module sub_7();
	    implement code
endmodule
