module sub_5();
	    implement code
endmodule
